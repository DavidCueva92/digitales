Library ieee;
Use ieee.std_logic_1164.all;
Use ieee.std_logic_unsigned.all;
Use IEEE.std_logic_arith.all;
Use work.mis_componentes.all;
---------------------------------------------------------------------------------------------------------
ENTITY REFLEJOS_HUMANOS IS
PORT(	START_P: 				In std_logic;
		BOTONERAS_P: 			In std_logic_vector(14 downto 0);
		RESET_P: 				In std_logic;
		CLOCK_FPGA: 		In std_logic;
		LEDS: 				Out std_logic_vector(14 downto 0);
		DEC_ACIERTOS:		Out std_logic_vector(6 downto 0);
		UNID_ACIERTOS:		Out std_logic_vector(6 downto 0);
		DEC_VELOCIDAD:		Out std_logic_vector(6 downto 0);
		UNID_VELOCIDAD:	Out std_logic_vector(6 downto 0));
END REFLEJOS_HUMANOS; 
---------------------------------------------------------------------------------------------------------
ARCHITECTURE estructural OF REFLEJOS_HUMANOS IS
-------------------------------------------------------------------------------------------------------------
TYPE ESTADO IS (T0, T1, T2, T3, T4, T5, T6, T7, T8);
SIGNAL Y: ESTADO;

SIGNAL START_N, RESET_N, START, RESET: std_logic;
SIGNAL BOTONERAS_N, BOTONERAS: std_logic_vector(14 downto 0);
SIGNAL RESET_CONT_1A15: std_logic;
SIGNAL EN_CONT_VECES, RESET_CONT_VECES, FIN_VECES: std_logic;
SIGNAL EN_REG, RESET_REG, DATA_CERO: std_logic;
SIGNAL NUM_1A15, VECES, NUM_LED: std_logic_vector(3 downto 0);
SIGNAL EN_CONT_15ds, RESET_CONT_15ds, IG_15ds: std_logic;
SIGNAL TIME_LED: std_logic_vector(3  downto 0);
SIGNAL SUMA_TIME, RESET_TIME: std_logic;
SIGNAL TIME_TOTAL: std_logic_vector(7 downto 0);
SIGNAL NUM_BOTONERA, NUM_TECLA: std_logic_vector(3 downto 0);
SIGNAL EN_REG_BOT, BOTON_PRESS, BOTON_OK: std_logic;
SIGNAL EN_CONT_ACIERTOS, RESET_CONT_ACIERTOS: std_logic;
SIGNAL ACIERTOS, DEC_BCD_ACIERT, UNID_BCD_ACIERT: std_logic_vector(3 downto 0);
SIGNAL EN_PROMEDIO, APAGAR: std_logic;
SIGNAL VELOCIDAD, DEC_BCD_VELOC, UNID_BCD_VELOC: std_logic_vector(3 downto 0);
SIGNAL SIN_USO_0, SIN_USO_1, SIN_USO_2: std_logic;
SIGNAL CLOCK_1MHz, CLOCK_100KHz, CLOCK_10KHz, CLOCK, CLOCK_100Hz, CLOCK_10Hz, CLOCK_1Hz: std_logic;
-------------------------------------------------------------------------------------------------------------
BEGIN
	MSS_TRANSICIONES: PROCESS(RESET, CLOCK)
	BEGIN
		IF RESET='1' THEN Y <= T0;
		ELSIF (CLOCK'EVENT AND CLOCK='1') THEN
			CASE Y IS
				WHEN T0 => IF START='0' THEN Y<=T0; ELSE Y<=T1; END IF;
				WHEN T1 => IF START='1' THEN Y<=T1; ELSE Y<=T2; END IF;
				WHEN T2 => IF FIN_VECES='1' THEN Y<=T3;
							  ELSIF DATA_CERO='0' THEN Y<=T4;
							  ELSE Y<=T2; END IF;
				WHEN T3 => IF START='0' THEN Y<=T3; ELSE Y<=T1; END IF;
				WHEN T4 => IF IG_15ds='1' THEN Y<=T5;
							  ELSIF BOTON_PRESS='1' THEN Y<=T7;
							  ELSE Y<=T4; END IF;
				WHEN T5 => Y<=T8;
				WHEN T6 => IF BOTON_OK='1' THEN Y<=T5; ELSE Y<=T8; END IF;
				WHEN T7 => IF BOTON_PRESS='0' THEN Y<=T6; ELSE Y<=T7; END IF;
				WHEN T8 => Y<=T2;
			END CASE;
		END IF;
	END PROCESS;
	
	MSS_SALIDAS: PROCESS(Y, START, FIN_VECES, DATA_CERO, IG_15ds, BOTON_PRESS, BOTON_OK)
	BEGIN
		RESET_CONT_1A15<='0'; RESET_TIME<='0'; RESET_CONT_VECES<='0'; RESET_REG<='0'; RESET_CONT_ACIERTOS<='0'; RESET_CONT_15ds<='0'; APAGAR<='0'; 
		EN_REG<='0'; EN_REG_BOT<='0'; EN_PROMEDIO<='0'; EN_CONT_15ds<='0'; SUMA_TIME<='0'; EN_CONT_ACIERTOS<='0'; EN_CONT_VECES<='0';
		CASE Y IS
			WHEN T0 =>  RESET_CONT_1A15<='1'; RESET_TIME<='1'; RESET_CONT_VECES<='1'; RESET_REG<='1'; RESET_CONT_ACIERTOS<='1'; RESET_CONT_15ds<='1'; APAGAR<='1'; 
			WHEN T1 =>  RESET_CONT_1A15<='1'; RESET_TIME<='1'; RESET_CONT_VECES<='1'; RESET_REG<='1'; RESET_CONT_ACIERTOS<='1'; RESET_CONT_15ds<='1'; APAGAR<='1'; 
			WHEN T2 =>  IF (FIN_VECES='0' AND DATA_CERO='1') THEN EN_REG<='1'; END IF;
			WHEN T3 =>  EN_PROMEDIO<='1';
			WHEN T4 =>  IF (IG_15ds='0' AND BOTON_PRESS='0') THEN EN_CONT_15ds<='1'; END IF;
			WHEN T5 =>  RESET_CONT_15ds<='1';
			WHEN T6 =>  IF BOTON_OK='1' THEN SUMA_TIME<='1'; EN_CONT_ACIERTOS<='1'; ELSE RESET_CONT_15ds<='1'; END IF;
			WHEN T7 =>  IF BOTON_PRESS='1' THEN EN_REG_BOT<='1'; END IF;
			WHEN T8 =>  RESET_REG<='1'; EN_CONT_VECES<='1';
		END CASE;
	END PROCESS;
	
	DIVISOR_FRECUENCIAS: CLOCK_DIV Port Map(CLOCK_FPGA, CLOCK_1MHz, CLOCK_100KHz, CLOCK_10KHz, CLOCK, CLOCK_100Hz, CLOCK_10Hz, CLOCK_1Hz);
	SIN_RIZADO_START: ANTIREBOTE Port Map (START_P, CLOCK_100Hz, START_N);
	SIN_RIZADO_RESET: ANTIREBOTE Port Map (RESET_P, CLOCK_100Hz, RESET_N);
	SIN_RIZADO_B1: ANTIREBOTE Port Map (BOTONERAS_P(0), CLOCK_100Hz, BOTONERAS_N(0));
	SIN_RIZADO_B2: ANTIREBOTE Port Map (BOTONERAS_P(1), CLOCK_100Hz, BOTONERAS_N(1));
	SIN_RIZADO_B3: ANTIREBOTE Port Map (BOTONERAS_P(2), CLOCK_100Hz, BOTONERAS_N(2));
	SIN_RIZADO_B4: ANTIREBOTE Port Map (BOTONERAS_P(3), CLOCK_100Hz, BOTONERAS_N(3));
	SIN_RIZADO_B5: ANTIREBOTE Port Map (BOTONERAS_P(4), CLOCK_100Hz, BOTONERAS_N(4));
	SIN_RIZADO_B6: ANTIREBOTE Port Map (BOTONERAS_P(5), CLOCK_100Hz, BOTONERAS_N(5));
	SIN_RIZADO_B7: ANTIREBOTE Port Map (BOTONERAS_P(6), CLOCK_100Hz, BOTONERAS_N(6));
	SIN_RIZADO_B8: ANTIREBOTE Port Map (BOTONERAS_P(7), CLOCK_100Hz, BOTONERAS_N(7));
	SIN_RIZADO_B9: ANTIREBOTE Port Map (BOTONERAS_P(8), CLOCK_100Hz, BOTONERAS_N(8));
	SIN_RIZADO_B10: ANTIREBOTE Port Map (BOTONERAS_P(9), CLOCK_100Hz, BOTONERAS_N(9));
	SIN_RIZADO_B11: ANTIREBOTE Port Map (BOTONERAS_P(10), CLOCK_100Hz, BOTONERAS_N(10));
	SIN_RIZADO_B12: ANTIREBOTE Port Map (BOTONERAS_P(11), CLOCK_100Hz, BOTONERAS_N(11));
	SIN_RIZADO_B13: ANTIREBOTE Port Map (BOTONERAS_P(12), CLOCK_100Hz, BOTONERAS_N(12));
	SIN_RIZADO_B14: ANTIREBOTE Port Map (BOTONERAS_P(13), CLOCK_100Hz, BOTONERAS_N(13));
	SIN_RIZADO_B15: ANTIREBOTE Port Map (BOTONERAS_P(14), CLOCK_100Hz, BOTONERAS_N(14));
	
	START <= NOT(START_N);
	RESET <= NOT(RESET_N);
	BOTONERAS(0) <= NOT(BOTONERAS_N(0));
	BOTONERAS(1) <= NOT(BOTONERAS_N(1));
	BOTONERAS(2) <= NOT(BOTONERAS_N(2));
	BOTONERAS(3) <= NOT(BOTONERAS_N(3));
	BOTONERAS(4) <= NOT(BOTONERAS_N(4));
	BOTONERAS(5) <= NOT(BOTONERAS_N(5));
	BOTONERAS(6) <= NOT(BOTONERAS_N(6));
	BOTONERAS(7) <= NOT(BOTONERAS_N(7));
	BOTONERAS(8) <= NOT(BOTONERAS_N(8));
	BOTONERAS(9) <= NOT(BOTONERAS_N(9));
	BOTONERAS(10) <= NOT(BOTONERAS_N(10));
	BOTONERAS(11) <= NOT(BOTONERAS_N(11));
	BOTONERAS(12) <= NOT(BOTONERAS_N(12));
	BOTONERAS(13) <= NOT(BOTONERAS_N(13));
	BOTONERAS(14) <= NOT(BOTONERAS_N(14));
	
	FIN_VECES <= (VECES(3) AND VECES(2) AND VECES(1) AND VECES(0));
	DATA_CERO <= NOT(NUM_LED(3) OR NUM_LED(2) OR NUM_LED(1) OR NUM_LED(0));
	BOTON_PRESS <= (BOTONERAS(14) OR BOTONERAS(13) OR BOTONERAS(12) OR BOTONERAS(11) OR BOTONERAS(10) OR BOTONERAS(9) OR BOTONERAS(8) OR BOTONERAS(7) OR BOTONERAS(6) OR BOTONERAS(5) OR BOTONERAS(4) OR BOTONERAS(3) OR BOTONERAS(2) OR BOTONERAS(1) OR BOTONERAS(0));
	IG_15ds <= (TIME_LED(3) AND TIME_LED(2) AND TIME_LED(1) AND TIME_LED(0));
	
	CONTADOR_UP_NUM1A15: CONTADOR_UP Port Map("0000", '1', '0', RESET_CONT_1A15, CLOCK_100Hz, NUM_1A15);
	REGISTRO_SOSTENIMIENTO_DIRECCION: REG_SOST Port Map(NUM_1A15, EN_REG, RESET_REG, CLOCK, NUM_LED);
	CONTADOR_UP_VECES: CONTADOR_UP Port Map("0000", EN_CONT_VECES, '0', RESET_CONT_VECES, CLOCK, VECES);
	DEMULTIPLEXADOR_LEDS: DEMUX_1TO16 Port Map('1', NUM_LED, SIN_USO_0, LEDS(0), LEDS(1), LEDS(2), LEDS(3), LEDS(4), LEDS(5), LEDS(6), LEDS(7), LEDS(8), LEDS(9), LEDS(10), LEDS(11), LEDS(12), LEDS(13), LEDS(14));
	CONTADOR_UP_TIME_LED: CONTADOR_UP Port Map("0000", EN_CONT_15ds, '0', RESET_CONT_15ds, CLOCK_10Hz, TIME_LED);
	SUMADOR_TIEMPO: SUMADOR_RETROALIMENTADO Port Map(TIME_LED, SUMA_TIME, '0', RESET_TIME, CLOCK, TIME_TOTAL);
	DECIMAL_A_BINARIO: DECODER_DECIMAL_BINARIO Port Map(BOTONERAS, NUM_BOTONERA);
	REGISTRO_SOSTENIMIENTO_BOTONERA: REG_SOST Port Map(NUM_BOTONERA, EN_REG_BOT, RESET_REG, CLOCK, NUM_TECLA);
	COMPARADOR_TECLA: COMPARADOR Port Map(NUM_LED, NUM_TECLA, SIN_USO_1, BOTON_OK, SIN_USO_2);
	CONTADOR_UP_ACIERTOS: CONTADOR_UP Port Map("0000", EN_CONT_ACIERTOS, '0', RESET_CONT_ACIERTOS, CLOCK, ACIERTOS);
	PROMEDIADOR: PROMEDIO Port Map(TIME_TOTAL, ACIERTOS, EN_PROMEDIO, VELOCIDAD);
	BINARIO_A_BCD_1: DECODER_BINARIO_BCD Port Map(VELOCIDAD, DEC_BCD_VELOC, UNID_BCD_VELOC);
	BINARIO_A_BCD_2: DECODER_BINARIO_BCD Port Map(ACIERTOS, DEC_BCD_ACIERT, UNID_BCD_ACIERT);
	VELOCIDAD_DECENAS: DECODER_7SEG Port Map(DEC_BCD_VELOC, APAGAR, DEC_VELOCIDAD);
	VELOCIDAD_UNIDADES: DECODER_7SEG Port Map(UNID_BCD_VELOC, APAGAR, UNID_VELOCIDAD);
	ACIERTOS_DECENAS: DECODER_7SEG Port Map(DEC_BCD_ACIERT, APAGAR, DEC_ACIERTOS);
	ACIERTOS_UNIDADES: DECODER_7SEG Port Map(UNID_BCD_ACIERT, APAGAR, UNID_ACIERTOS);
	
END estructural;


	